module reset( input clk,
              input rst_l_in,
              input rst_l_out)
);
